//  Module: or_module
//

module or_module
    (
        input logic a,
        input logic b,
        output logic y
    );

    assign y = a || b;
endmodule: or_module
